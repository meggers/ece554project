module ID_Unit(clk, rst);

//////////////////////////INPUTS/////////////////////////////

/////////////////////////END INPUTS///////////////////////////

//////////////////////////OUTPUTS/////////////////////////////

////////////////////////END OUTPUTS///////////////////////////
                
endmodule
