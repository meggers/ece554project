library verilog;
use verilog.vl_types.all;
entity BasicOp_tb is
end BasicOp_tb;
