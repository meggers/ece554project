// Author: Graham Nygard, Robert Wagner

module IDEX_reg(clk);

//INPUTS/////////////////////////////

//OUTPUTS/////////////////////////////

endmodule
