module EX_Unit(clk);

//////////////////////////INPUTS/////////////////////////////

/////////////////////////END INPUTS///////////////////////////

//////////////////////////OUTPUTS/////////////////////////////

////////////////////////END OUTPUTS///////////////////////////

endmodule
