library verilog;
use verilog.vl_types.all;
entity Control_tb is
end Control_tb;
