library verilog;
use verilog.vl_types.all;
entity Full_processor_v_unit is
end Full_processor_v_unit;
