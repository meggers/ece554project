library verilog;
use verilog.vl_types.all;
entity Loop_tb is
end Loop_tb;
