library verilog;
use verilog.vl_types.all;
entity Full_processor_tb is
end Full_processor_tb;
