library verilog;
use verilog.vl_types.all;
entity DataDependence_tb is
end DataDependence_tb;
