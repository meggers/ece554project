module reg_file(p0, p1, re0, re1, p0_addr, p1_addr, dst_addr, dst, WE, clk,
                  bus_out0, bus_out1, bus_out2, bus_out3, bus_out4, 
                  bus_out5, bus_out6, bus_out7, bus_out8, bus_out9,
                  bus_out10, bus_out11, bus_out12, bus_out13, bus_out14,
                  bus_out15);
   output [15:0] p0, p1; 
   input [15:0] dst; 
   input [3:0] p0_addr, p1_addr, dst_addr;
   input WE, clk, re0, re1;
   
   localparam R0 = 4'h0;
   localparam R1 = 4'h1;
   localparam R2 = 4'h2;
   localparam R3 = 4'h3; 
   localparam R4 = 4'h4; 
   localparam R5 = 4'h5; 
   localparam R6 = 4'h6; 
   localparam R7 = 4'h7; 
   localparam R8 = 4'h8; 
   localparam R9 = 4'h9; 
   localparam R10 = 4'hA; 
   localparam R11 = 4'hB; 
   localparam R12 = 4'hC; 
   localparam R13 = 4'hD; 
   localparam R14 = 4'hE; 
   localparam R15 = 4'hF; 
   
   
   //input write signals to registers
   reg [15:0] rw;
                  
   //outputs of registers
   output [15:0] bus_out0, bus_out1, bus_out2, bus_out3, bus_out4, 
                  bus_out5, bus_out6, bus_out7, bus_out8, bus_out9,
                  bus_out10, bus_out11, bus_out12, bus_out13, bus_out14,
                  bus_out15;
   
   
   Reg16 r0(.bus_out(bus_out0), .regWrite(rw[0]), .bus_in(dst), .clk(clk));
   Reg16 r1(.bus_out(bus_out1), .regWrite(rw[1]), .bus_in(dst), .clk(clk)); 
   Reg16 r2(.bus_out(bus_out2), .regWrite(rw[2]), .bus_in(dst), .clk(clk)); 
   Reg16 r3(.bus_out(bus_out3), .regWrite(rw[3]), .bus_in(dst), .clk(clk)); 
   Reg16 r4(.bus_out(bus_out4), .regWrite(rw[4]), .bus_in(dst), .clk(clk)); 
   Reg16 r5(.bus_out(bus_out5), .regWrite(rw[5]), .bus_in(dst), .clk(clk)); 
   Reg16 r6(.bus_out(bus_out6), .regWrite(rw[6]), .bus_in(dst), .clk(clk));  
   Reg16 r7(.bus_out(bus_out7), .regWrite(rw[7]), .bus_in(dst), .clk(clk));
   Reg16 r8(.bus_out(bus_out8), .regWrite(rw[8]), .bus_in(dst), .clk(clk)); 
   Reg16 r9(.bus_out(bus_out9), .regWrite(rw[9]), .bus_in(dst), .clk(clk)); 
   Reg16 r10(.bus_out(bus_out10), .regWrite(rw[10]), .bus_in(dst), .clk(clk)); 
   Reg16 r11(.bus_out(bus_out11), .regWrite(rw[11]), .bus_in(dst), .clk(clk));
   Reg16 r12(.bus_out(bus_out12), .regWrite(rw[12]), .bus_in(dst), .clk(clk)); 
   Reg16 r13(.bus_out(bus_out13), .regWrite(rw[13]), .bus_in(dst), .clk(clk));
   Reg16 r14(.bus_out(bus_out14), .regWrite(rw[14]), .bus_in(dst), .clk(clk)); 
   Reg16 r15(.bus_out(bus_out15), .regWrite(rw[15]), .bus_in(dst), .clk(clk));
   
   assign p0 = ((p0_addr == R0) && (re0)) ? bus_out0:
                 ((p0_addr == R1) && (re0)) ? bus_out1:
                 ((p0_addr == R2) && (re0)) ? bus_out2:
                 ((p0_addr == R3) && (re0)) ? bus_out3:
                 ((p0_addr == R4) && (re0)) ? bus_out4:
                 ((p0_addr == R5) && (re0)) ? bus_out5:
                 ((p0_addr == R6) && (re0)) ? bus_out6:
                 ((p0_addr == R7) && (re0)) ? bus_out7:
                 ((p0_addr == R8) && (re0)) ? bus_out8:
                 ((p0_addr == R9) && (re0)) ? bus_out9:
                 ((p0_addr == R10) && (re0)) ? bus_out10:
                 ((p0_addr == R11) && (re0)) ? bus_out11:
                 ((p0_addr == R12) && (re0)) ? bus_out12:
                 ((p0_addr == R13) && (re0)) ? bus_out13:
                 ((p0_addr == R14) && (re0)) ? bus_out14:
                 ((p0_addr == R15) && (re0)) ? bus_out15:
					    16'hxxxx;
   
   assign p1 = ((p1_addr == R0) && (re1)) ? bus_out0:
                 ((p1_addr == R1) && (re1)) ? bus_out1:
                 ((p1_addr == R2) && (re1)) ? bus_out2:
                 ((p1_addr == R3) && (re1)) ? bus_out3:
                 ((p1_addr == R4) && (re1)) ? bus_out4:
                 ((p1_addr == R5) && (re1)) ? bus_out5:
                 ((p1_addr == R6) && (re1)) ? bus_out6:
                 ((p1_addr == R7) && (re1)) ? bus_out7:
                 ((p1_addr == R8) && (re1)) ? bus_out8:
                 ((p1_addr == R9) && (re1)) ? bus_out9:
                 ((p1_addr == R10) && (re1)) ? bus_out10:
                 ((p1_addr == R11) && (re1)) ? bus_out11:
                 ((p1_addr == R12) && (re1)) ? bus_out12:
                 ((p1_addr == R13) && (re1)) ? bus_out13:
                 ((p1_addr == R14) && (re1)) ? bus_out14:
                 ((p1_addr == R15) && (re1)) ? bus_out15:
					    16'hxxxx;
                                  
    always @(dst_addr, WE) begin
        if(WE) 
           case (dst_addr)
               R0: rw = 16'h0001;
               R1: rw = 16'h0002;
               R2: rw = 16'h0004;
               R3: rw = 16'h0008;
               R4: rw = 16'h0010;
               R5: rw = 16'h0020;
               R6: rw = 16'h0040;
               R7: rw = 16'h0080;
               R8: rw = 16'h0100;
               R9: rw = 16'h0200;
               R10: rw = 16'h0400;
               R11: rw = 16'h0800;
               R12: rw = 16'h1000;
               R13: rw = 16'h2000;
               R14: rw = 16'h4000;
               R15: rw = 16'h8000;
          endcase 
       else
          rw = 16'h0000;

   end 
   
endmodule 
       
       
       