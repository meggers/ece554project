library verilog;
use verilog.vl_types.all;
entity datapath is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        instr           : in     vl_logic_vector(15 downto 0);
        p0_addr         : out    vl_logic_vector(3 downto 0);
        p1_addr         : out    vl_logic_vector(3 downto 0);
        p0              : in     vl_logic_vector(15 downto 0);
        p1              : in     vl_logic_vector(15 downto 0);
        dst             : out    vl_logic_vector(15 downto 0);
        dst_addr        : out    vl_logic_vector(3 downto 0);
        WE              : out    vl_logic;
        hlt             : out    vl_logic;
        op_ALU          : out    vl_logic_vector(3 downto 0);
        ALU_mux         : in     vl_logic_vector(3 downto 0);
        reg0_addr_cntrl : in     vl_logic_vector(2 downto 0);
        reg1_addr_cntrl : in     vl_logic_vector(2 downto 0);
        load_LH_sel     : in     vl_logic;
        dst_sel         : in     vl_logic_vector(2 downto 0);
        dst_addr_sel    : in     vl_logic_vector(2 downto 0);
        WE_cntrl        : in     vl_logic;
        \WE_DM\         : in     vl_logic;
        \RE_DM\         : in     vl_logic;
        we_dm           : out    vl_logic;
        re_dm           : out    vl_logic;
        PC_mux          : in     vl_logic_vector(1 downto 0);
        RE_0            : in     vl_logic;
        RE_1            : in     vl_logic;
        IFID            : out    vl_logic_vector(15 downto 0);
        Bad_Instr_CNTRL : in     vl_logic;
        Bad_Instr_IDEX  : out    vl_logic;
        b_true          : in     vl_logic;
        PC_mux_RET      : in     vl_logic;
        Bad_Instr_RET   : in     vl_logic;
        Bad_Instr_RET_IDEX: out    vl_logic;
        Bad_Instr_RET_EXMEM: out    vl_logic;
        Bad_Instr_RET_IFID: out    vl_logic;
        call_ret_hold_bad: out    vl_logic;
        ALU_out         : in     vl_logic_vector(15 downto 0);
        ALU_in1         : out    vl_logic_vector(15 downto 0);
        ALU_in2         : out    vl_logic_vector(15 downto 0);
        addr_DM         : out    vl_logic_vector(15 downto 0);
        addr_DM_mux     : in     vl_logic_vector(3 downto 0);
        rd_DM           : in     vl_logic_vector(15 downto 0);
        wd_dm           : out    vl_logic_vector(15 downto 0);
        PC              : out    vl_logic_vector(15 downto 0);
        No_Op_IFID      : in     vl_logic;
        No_Op_IDEX      : out    vl_logic;
        rd_rt_addr_IDEX : out    vl_logic_vector(3 downto 0);
        rd_rt_addr_EXMEM: out    vl_logic_vector(3 downto 0);
        rd_rt_addr_MEMWB: out    vl_logic_vector(3 downto 0);
        rd_rt_addr_WB   : out    vl_logic_vector(3 downto 0);
        pc_stop_icache_mem: in     vl_logic;
        we_icache       : in     vl_logic;
        dataforward_EXMEM_P0_ff: in     vl_logic;
        dataforward_EXMEM_P1_ff: in     vl_logic;
        dataforward_MEMWB_P0_ff: in     vl_logic;
        dataforward_MEMWB_P1_ff: in     vl_logic;
        dataforward_WB_P0_ff: in     vl_logic;
        dataforward_WB_P1_ff: in     vl_logic
    );
end datapath;
