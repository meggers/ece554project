module IF_Unit(clk, rst, data_hazard, instruction);

//////////////////////////INPUTS/////////////////////////////

/////////////////////////END INPUTS///////////////////////////

//////////////////////////OUTPUTS/////////////////////////////

////////////////////////END OUTPUTS///////////////////////////

endmodule
