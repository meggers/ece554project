library verilog;
use verilog.vl_types.all;
entity control is
    port(
        IFID            : in     vl_logic_vector(15 downto 0);
        rst             : in     vl_logic;
        clk             : in     vl_logic;
        WE              : out    vl_logic;
        ALU_mux         : out    vl_logic_vector(3 downto 0);
        reg0_addr_cntrl : out    vl_logic_vector(2 downto 0);
        reg1_addr_cntrl : out    vl_logic_vector(2 downto 0);
        RE_0            : out    vl_logic;
        RE_1            : out    vl_logic;
        N               : in     vl_logic;
        Z               : in     vl_logic;
        V               : in     vl_logic;
        load_LH_sel     : out    vl_logic;
        dst_sel         : out    vl_logic_vector(2 downto 0);
        dst_addr_sel    : out    vl_logic_vector(2 downto 0);
        WE_DM           : out    vl_logic;
        RE_DM           : out    vl_logic;
        addr_DM_mux     : out    vl_logic_vector(3 downto 0);
        rd_en_IM        : out    vl_logic;
        PC_mux          : out    vl_logic_vector(1 downto 0);
        No_Op_IFID      : out    vl_logic;
        p0_addr         : in     vl_logic_vector(3 downto 0);
        p1_addr         : in     vl_logic_vector(3 downto 0);
        dst_addr_IDEX   : in     vl_logic_vector(3 downto 0);
        dst_addr_EXMEM  : in     vl_logic_vector(3 downto 0);
        dst_addr_MEMWB  : in     vl_logic_vector(3 downto 0);
        dst_addr_WB     : in     vl_logic_vector(3 downto 0);
        No_Op_IDEX      : in     vl_logic;
        Bad_Instr       : out    vl_logic;
        Bad_Instr_IDEX  : in     vl_logic;
        b_true          : out    vl_logic;
        PC_mux_RET      : out    vl_logic;
        Bad_Instr_RET   : out    vl_logic;
        Bad_Instr_RET_IDEX: in     vl_logic;
        Bad_Instr_RET_EXMEM: in     vl_logic;
        Bad_Instr_RET_IFID: in     vl_logic;
        call_ret_hold_bad: in     vl_logic;
        no_op_icache    : in     vl_logic;
        N_ff            : out    vl_logic;
        Z_ff            : out    vl_logic;
        V_ff            : out    vl_logic;
        instr_go        : in     vl_logic;
        dataforward_EXMEM_P0_ff: out    vl_logic;
        dataforward_EXMEM_P1_ff: out    vl_logic;
        dataforward_MEMWB_P0_ff: out    vl_logic;
        dataforward_MEMWB_P1_ff: out    vl_logic;
        dataforward_WB_P0_ff: out    vl_logic;
        dataforward_WB_P1_ff: out    vl_logic
    );
end control;
