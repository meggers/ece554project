library verilog;
use verilog.vl_types.all;
entity Branch_tb is
end Branch_tb;
