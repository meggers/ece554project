// Author: Graham Nygard, Robert Wagner

module IDEX_reg(clk);

//////////////////////////INPUTS/////////////////////////////

/////////////////////////END INPUTS///////////////////////////

//////////////////////////OUTPUTS/////////////////////////////

////////////////////////END OUTPUTS///////////////////////////

endmodule
