module WB_Unit();

///////////////////////////INPUTS/////////////////////////////

/////////////////////////END INPUTS///////////////////////////

//////////////////////////OUTPUTS/////////////////////////////

////////////////////////END OUTPUTS///////////////////////////

endmodule
