library verilog;
use verilog.vl_types.all;
entity LwStall_tb is
end LwStall_tb;
